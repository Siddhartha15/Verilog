module encoder
	
endmodule
